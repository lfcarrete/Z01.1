-- Elementos de Sistemas
-- by Luciano Soares
-- HalfAdder.vhd

-- Implementa Half Adder

Library ieee;
use ieee.std_logic_1164.all;

entity HalfAdder is
	port(
		a,b:         in STD_LOGIC;   -- entradas
		soma,vaium: out STD_LOGIC   -- sum e carry
	);
end entity;

architecture rtl of HalfAdder is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.

begin
<<<<<<< HEAD
  -- Implementação vem aqui!
  soma <= a xor b;
=======
  
  soma <= (a and not(b)) or (not(a) and b);

>>>>>>> ULAupgrade
  vaium <= a and b;

end architecture;
